magic
tech sky130A
timestamp 1614729275
<< nwell >>
rect -150 90 510 485
<< nmos >>
rect -35 -90 -20 10
rect 110 -90 125 10
rect 255 -90 315 10
rect 445 -90 460 10
rect 110 -340 125 -240
rect 255 -340 315 -240
rect 445 -340 460 -240
<< pmos >>
rect -80 365 -20 465
rect 110 365 125 465
rect 255 365 270 465
rect 320 365 335 465
rect -80 110 -20 210
rect 110 110 125 210
rect 320 110 335 210
<< ndiff >>
rect -85 -10 -35 10
rect -85 -70 -70 -10
rect -50 -70 -35 -10
rect -85 -90 -35 -70
rect -20 -10 30 10
rect -20 -70 -5 -10
rect 15 -70 30 -10
rect -20 -90 30 -70
rect 60 -10 110 10
rect 60 -70 75 -10
rect 95 -70 110 -10
rect 60 -90 110 -70
rect 125 -10 175 10
rect 125 -70 140 -10
rect 160 -70 175 -10
rect 125 -90 175 -70
rect 205 -10 255 10
rect 205 -70 220 -10
rect 240 -70 255 -10
rect 205 -90 255 -70
rect 315 -10 365 10
rect 315 -70 330 -10
rect 350 -70 365 -10
rect 315 -90 365 -70
rect 395 -10 445 10
rect 395 -70 410 -10
rect 430 -70 445 -10
rect 395 -90 445 -70
rect 460 -10 510 10
rect 460 -70 475 -10
rect 495 -70 510 -10
rect 460 -90 510 -70
rect 60 -260 110 -240
rect 60 -320 75 -260
rect 95 -320 110 -260
rect 60 -340 110 -320
rect 125 -260 175 -240
rect 125 -320 140 -260
rect 160 -320 175 -260
rect 125 -340 175 -320
rect 205 -260 255 -240
rect 205 -320 220 -260
rect 240 -320 255 -260
rect 205 -340 255 -320
rect 315 -260 365 -240
rect 315 -320 330 -260
rect 350 -320 365 -260
rect 315 -340 365 -320
rect 395 -260 445 -240
rect 395 -320 410 -260
rect 430 -320 445 -260
rect 395 -340 445 -320
rect 460 -260 510 -240
rect 460 -320 475 -260
rect 495 -320 510 -260
rect 460 -340 510 -320
<< pdiff >>
rect -130 445 -80 465
rect -130 385 -115 445
rect -95 385 -80 445
rect -130 365 -80 385
rect -20 445 30 465
rect -20 385 -5 445
rect 15 385 30 445
rect -20 365 30 385
rect 60 445 110 465
rect 60 385 75 445
rect 95 385 110 445
rect 60 365 110 385
rect 125 445 175 465
rect 125 385 140 445
rect 160 385 175 445
rect 125 365 175 385
rect 205 445 255 465
rect 205 385 220 445
rect 240 385 255 445
rect 205 365 255 385
rect 270 445 320 465
rect 270 385 285 445
rect 305 385 320 445
rect 270 365 320 385
rect 335 445 385 465
rect 335 385 350 445
rect 370 385 385 445
rect 335 365 385 385
rect -130 190 -80 210
rect -130 130 -115 190
rect -95 130 -80 190
rect -130 110 -80 130
rect -20 190 30 210
rect -20 130 -5 190
rect 15 130 30 190
rect -20 110 30 130
rect 60 190 110 210
rect 60 130 75 190
rect 95 130 110 190
rect 60 110 110 130
rect 125 190 175 210
rect 125 130 140 190
rect 160 130 175 190
rect 125 110 175 130
rect 270 190 320 210
rect 270 130 285 190
rect 305 130 320 190
rect 270 110 320 130
rect 335 190 385 210
rect 335 130 350 190
rect 370 130 385 190
rect 335 110 385 130
<< ndiffc >>
rect -70 -70 -50 -10
rect -5 -70 15 -10
rect 75 -70 95 -10
rect 140 -70 160 -10
rect 220 -70 240 -10
rect 330 -70 350 -10
rect 410 -70 430 -10
rect 475 -70 495 -10
rect 75 -320 95 -260
rect 140 -320 160 -260
rect 220 -320 240 -260
rect 330 -320 350 -260
rect 410 -320 430 -260
rect 475 -320 495 -260
<< pdiffc >>
rect -115 385 -95 445
rect -5 385 15 445
rect 75 385 95 445
rect 140 385 160 445
rect 220 385 240 445
rect 285 385 305 445
rect 350 385 370 445
rect -115 130 -95 190
rect -5 130 15 190
rect 75 130 95 190
rect 140 130 160 190
rect 285 130 305 190
rect 350 130 370 190
<< psubdiff >>
rect -135 -10 -85 10
rect -135 -70 -120 -10
rect -100 -70 -85 -10
rect -135 -90 -85 -70
<< nsubdiff >>
rect 415 190 465 210
rect 415 130 430 190
rect 450 130 465 190
rect 415 110 465 130
<< psubdiffcont >>
rect -120 -70 -100 -10
<< nsubdiffcont >>
rect 430 130 450 190
<< poly >>
rect -80 465 -20 480
rect 110 465 125 480
rect 255 465 270 480
rect 320 465 335 480
rect -80 350 -20 365
rect -80 225 -65 350
rect 5 340 45 350
rect 5 320 15 340
rect 35 320 45 340
rect 5 310 45 320
rect 110 310 125 365
rect 170 340 210 350
rect 170 320 180 340
rect 200 320 210 340
rect 170 310 210 320
rect 30 240 45 310
rect 105 300 145 310
rect 105 280 115 300
rect 135 280 145 300
rect 105 270 145 280
rect 170 240 185 310
rect 30 225 185 240
rect 255 235 270 365
rect 320 310 335 365
rect 380 340 420 350
rect 380 320 390 340
rect 410 320 420 340
rect 380 310 420 320
rect 315 300 355 310
rect 315 280 325 300
rect 345 280 355 300
rect 315 270 355 280
rect 380 240 395 310
rect -80 210 -20 225
rect 110 210 125 225
rect 230 220 270 235
rect 320 225 395 240
rect -80 95 -20 110
rect -35 10 -20 95
rect 110 40 125 110
rect 230 100 245 220
rect 320 210 335 225
rect 230 85 270 100
rect 180 55 220 65
rect 180 40 190 55
rect 110 35 190 40
rect 210 35 220 55
rect 110 25 220 35
rect 255 25 270 85
rect 320 65 335 110
rect 445 85 485 95
rect 445 65 455 85
rect 475 65 485 85
rect 320 50 355 65
rect 340 40 355 50
rect 445 55 485 65
rect 445 40 460 55
rect 340 25 460 40
rect 110 10 125 25
rect 255 10 315 25
rect 445 10 460 25
rect -35 -105 -20 -90
rect 110 -100 125 -90
rect -75 -115 -20 -105
rect -75 -135 -65 -115
rect -45 -120 -20 -115
rect 25 -115 65 -105
rect -45 -135 -35 -120
rect -75 -145 -35 -135
rect 25 -135 35 -115
rect 55 -135 65 -115
rect 25 -145 65 -135
rect 110 -110 230 -100
rect 110 -115 200 -110
rect 110 -145 125 -115
rect 190 -130 200 -115
rect 220 -130 230 -110
rect 190 -140 230 -130
rect 255 -105 315 -90
rect 50 -210 65 -145
rect 90 -155 130 -145
rect 90 -175 100 -155
rect 120 -175 130 -155
rect 90 -185 130 -175
rect 190 -195 230 -185
rect 190 -210 200 -195
rect 50 -215 200 -210
rect 220 -215 230 -195
rect 50 -225 230 -215
rect 255 -225 270 -105
rect 360 -115 400 -105
rect 360 -135 370 -115
rect 390 -135 400 -115
rect 360 -145 400 -135
rect 445 -145 460 -90
rect 385 -210 400 -145
rect 425 -155 465 -145
rect 425 -175 435 -155
rect 455 -175 465 -155
rect 425 -185 465 -175
rect 385 -225 460 -210
rect 110 -240 125 -225
rect 255 -240 315 -225
rect 445 -240 460 -225
rect 110 -355 125 -340
rect 255 -355 315 -340
rect 445 -355 460 -340
rect 255 -365 295 -355
rect 255 -385 265 -365
rect 285 -385 295 -365
rect 255 -395 295 -385
<< polycont >>
rect 15 320 35 340
rect 180 320 200 340
rect 115 280 135 300
rect 390 320 410 340
rect 325 280 345 300
rect 190 35 210 55
rect 455 65 475 85
rect -65 -135 -45 -115
rect 35 -135 55 -115
rect 200 -130 220 -110
rect 100 -175 120 -155
rect 200 -215 220 -195
rect 370 -135 390 -115
rect 435 -175 455 -155
rect 265 -385 285 -365
<< locali >>
rect -125 445 -85 460
rect -125 390 -115 445
rect -150 385 -115 390
rect -95 385 -85 445
rect -150 370 -85 385
rect -15 445 25 460
rect -15 385 -5 445
rect 15 385 25 445
rect -15 370 25 385
rect 5 350 25 370
rect 65 445 105 460
rect 65 385 75 445
rect 95 385 105 445
rect 65 370 105 385
rect 130 445 170 460
rect 130 385 140 445
rect 160 385 170 445
rect 130 370 170 385
rect 210 445 250 460
rect 210 385 220 445
rect 240 385 250 445
rect 210 370 250 385
rect 275 445 315 460
rect 275 385 285 445
rect 305 385 315 445
rect 275 370 315 385
rect 340 445 380 460
rect 340 385 350 445
rect 370 385 380 445
rect 340 370 380 385
rect 5 340 45 350
rect 5 320 15 340
rect 35 320 45 340
rect 5 310 45 320
rect 65 205 85 370
rect 150 350 170 370
rect 150 340 210 350
rect 150 330 180 340
rect 170 320 180 330
rect 200 320 210 340
rect 170 310 210 320
rect 105 300 145 310
rect 105 280 115 300
rect 135 290 145 300
rect 135 280 170 290
rect 105 270 170 280
rect 150 205 170 270
rect -125 190 -85 205
rect -125 130 -115 190
rect -95 130 -85 190
rect -125 115 -85 130
rect -15 190 25 205
rect -15 130 -5 190
rect 15 130 25 190
rect -15 115 25 130
rect 65 190 105 205
rect 65 130 75 190
rect 95 130 105 190
rect 65 115 105 130
rect 130 190 170 205
rect 130 130 140 190
rect 160 130 170 190
rect 130 115 170 130
rect 275 205 295 370
rect 360 350 380 370
rect 450 370 510 390
rect 360 340 420 350
rect 360 330 390 340
rect 380 320 390 330
rect 410 320 420 340
rect 380 310 420 320
rect 315 300 355 310
rect 315 280 325 300
rect 345 290 355 300
rect 450 290 470 370
rect 345 280 470 290
rect 315 270 470 280
rect 360 205 380 270
rect 275 190 315 205
rect 275 130 285 190
rect 305 130 315 190
rect 275 115 315 130
rect 340 190 380 205
rect 340 130 350 190
rect 370 130 380 190
rect 340 115 380 130
rect 420 190 460 205
rect 420 130 430 190
rect 450 130 460 190
rect 420 115 460 130
rect -125 95 -105 115
rect -150 75 -105 95
rect 5 85 25 115
rect 130 85 150 115
rect 5 65 150 85
rect 65 5 85 65
rect 180 55 220 65
rect 180 35 190 55
rect 210 45 220 55
rect 210 35 230 45
rect 180 25 230 35
rect 210 5 230 25
rect 340 5 360 115
rect 445 85 510 95
rect 445 65 455 85
rect 475 75 510 85
rect 475 65 485 75
rect 445 55 485 65
rect -130 -10 -40 5
rect -130 -70 -120 -10
rect -100 -70 -70 -10
rect -50 -70 -40 -10
rect -130 -85 -40 -70
rect -15 -10 25 5
rect -15 -70 -5 -10
rect 15 -70 25 -10
rect -15 -85 25 -70
rect 65 -10 105 5
rect 65 -70 75 -10
rect 95 -70 105 -10
rect 65 -85 105 -70
rect 130 -10 170 5
rect 130 -70 140 -10
rect 160 -70 170 -10
rect 130 -85 170 -70
rect -75 -115 -35 -105
rect -75 -135 -65 -115
rect -45 -135 -35 -115
rect -75 -145 -35 -135
rect -55 -395 -35 -145
rect -15 -355 5 -85
rect 65 -105 85 -85
rect 25 -115 85 -105
rect 25 -135 35 -115
rect 55 -125 85 -115
rect 55 -135 65 -125
rect 25 -145 65 -135
rect 90 -155 130 -145
rect 90 -165 100 -155
rect 65 -175 100 -165
rect 120 -175 130 -155
rect 65 -185 130 -175
rect 65 -245 85 -185
rect 150 -245 170 -85
rect 210 -10 250 5
rect 210 -70 220 -10
rect 240 -70 250 -10
rect 210 -85 250 -70
rect 320 -10 440 5
rect 320 -70 330 -10
rect 350 -15 410 -10
rect 350 -70 360 -15
rect 320 -85 360 -70
rect 400 -70 410 -15
rect 430 -70 440 -10
rect 400 -85 440 -70
rect 465 -10 505 5
rect 465 -70 475 -10
rect 495 -70 505 -10
rect 465 -85 505 -70
rect 210 -100 230 -85
rect 190 -110 230 -100
rect 400 -105 420 -85
rect 190 -130 200 -110
rect 220 -130 230 -110
rect 190 -140 230 -130
rect 360 -115 420 -105
rect 360 -135 370 -115
rect 390 -125 420 -115
rect 390 -135 400 -125
rect 360 -145 400 -135
rect 425 -155 465 -145
rect 425 -165 435 -155
rect 400 -175 435 -165
rect 455 -175 465 -155
rect 400 -185 465 -175
rect 190 -195 230 -185
rect 190 -215 200 -195
rect 220 -215 230 -195
rect 190 -225 230 -215
rect 65 -260 105 -245
rect 65 -320 75 -260
rect 95 -320 105 -260
rect 65 -335 105 -320
rect 130 -260 170 -245
rect 130 -320 140 -260
rect 160 -320 170 -260
rect 130 -335 170 -320
rect 210 -245 230 -225
rect 400 -245 420 -185
rect 485 -245 505 -85
rect 210 -260 250 -245
rect 210 -320 220 -260
rect 240 -320 250 -260
rect 210 -335 250 -320
rect 320 -260 440 -245
rect 320 -320 330 -260
rect 350 -265 410 -260
rect 350 -320 360 -265
rect 320 -335 360 -320
rect 400 -320 410 -265
rect 430 -320 440 -260
rect 400 -335 440 -320
rect 465 -260 505 -245
rect 465 -320 475 -260
rect 495 -320 505 -260
rect 465 -335 505 -320
rect 130 -355 150 -335
rect -15 -375 150 -355
rect 255 -365 295 -355
rect 255 -385 265 -365
rect 285 -385 295 -365
rect 255 -395 295 -385
rect -150 -415 510 -395
<< viali >>
rect 75 385 95 445
rect 220 385 240 445
rect 75 130 95 190
rect 430 130 450 190
rect -120 -70 -100 -10
rect -70 -70 -50 -10
rect 475 -70 495 -10
rect 475 -320 495 -260
<< metal1 >>
rect -150 445 510 460
rect -150 385 75 445
rect 95 385 220 445
rect 240 385 510 445
rect -150 370 510 385
rect 65 190 105 370
rect 65 130 75 190
rect 95 130 105 190
rect 65 115 105 130
rect 420 190 460 370
rect 420 130 430 190
rect 450 130 460 190
rect 420 115 460 130
rect -150 -10 510 5
rect -150 -70 -120 -10
rect -100 -70 -70 -10
rect -50 -70 475 -10
rect 495 -70 510 -10
rect -150 -85 510 -70
rect 465 -260 505 -85
rect 465 -320 475 -260
rect 495 -320 505 -260
rect 465 -335 505 -320
<< labels >>
rlabel metal1 -150 415 -150 415 7 VP
port 1 w
rlabel locali -150 380 -150 380 7 D
port 5 w
rlabel locali -150 85 -150 85 7 Dn
port 6 w
rlabel locali -150 -405 -150 -405 7 CLK
port 3 w
rlabel metal1 -150 -40 -150 -40 7 VN
port 2 w
rlabel locali 510 380 510 380 3 Q
port 7 e
rlabel locali 510 85 510 85 3 Qn
port 8 e
<< end >>
